`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////

// inout f; to declare if it is an input and out 
// module myand (input a,b, 
//               output c);
module myand(a,b,c);
    input a,b;
    output c;
    
    and g1(c,a,b);
    
endmodule
